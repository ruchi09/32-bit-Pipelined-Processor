module piplinedprefix_tb();

reg [31:0]a,b;
reg c,clk;

wire [31:0]s;
wire cout;

prefix32 p(a,b,c,cout,s,clk);
initial
begin
clk=0;
end

always
begin
#1
clk=~clk;
end

initial

begin

#2
a=32'd23;
b=32'd11;
c=1;

/*
#2
a=32'd99;
b=32'd100;
c=1;


#2
a=32'd55;
b=32'd44;
c=1;


#2
a=32'd9;
b=32'd1;
c=0;

#2
a=32'b00000000000000000000000000000100;
b=32'b00000000000000000000000001000000;
c=1;


#2
a=32'b00000000000000000000000000000000;
b=32'b00000000000000000000000011111111;
c=1;


#2
a=32'b00000000000000000000000001111100;
b=32'b00000000000000000000000001000000;
c=1;
/*
#2
a=32'b00000000111100001111000000000000;
b=32'b00001111000000000000111100000000;
c=0;

#2
a=32'b11110000111100001111000011110000;
b=32'b00001111000011110000111100001111;
c=0;

#2
a=32'b11110000111100001111000011110000;
b=32'b00001111000011110000111100001111;
c=1;


*/
end



always 
begin
#23 $finish;
end 


initial
begin
$monitor($time,"\ns=%b  cout=%d  a=%d  b=%d  c=%d \n",s,cout,a,b,c );
end
endmodule

module mul_tb();

reg [31:0]x,y;
reg clk;

wire [63:0]s;
wire cout,cout1;

mul mul32(x,y,s,cout,clk,cout1);
initial
begin
clk=0;
end

always
begin
#1
clk=~clk;
end

initial

begin

#2
y=32'd1111;
x=32'd0;

/*
#2
y=32'd11111;
x=32'd10;


#2
y=32'd111;
x=32'd111;


#2
y=32'd22;
x=32'd22;


#2
y=32'd505000;
x=32'd100;

/*
#2
y=32'b00000000000000000000000000111111;
x=32'b100000;


#2
y=32'b00000000000000000000000000111111;
x=32'b1000000;



#2
y=32'b00000000000000000000000000111111;
x=32'b10000000;

#2
y=32'b00000000000000000000000000111111;
x=32'b100000000;

#2
y=32'b00000000000000000000000000111111;
x=32'b1000000000;
    
#2
y=32'b00000000000000000000000000111111;
x=32'b10000000000;


#2
y=32'b00000000000000000000000000111111;
x=32'b100000000000;


#2
y=32'b00000000000000000000000000111111;
x=32'b1000000000000;

#2
y=32'b00000000000000000000000000111111;
x=32'b10000000000000;


#2
y=32'b00000000000000000000000000111111;
x=32'b100000000000000;

#2
y=32'b00000000000000000000000000111111;
x=32'b1000000000000000;


#2
y=32'b00000000000000000000000000111111;
x=32'b10000000000000000;


#2
y=32'b00000000000000000000000000111111;
x=32'b10000000000000000000000000000;

#2
y=32'b00000000000000000000000000111111;
x=32'b100000000000000000000000000000;

#2
y=32'b00000000000000000000000000111111;
x=32'b1000000000000000000000000000000;

#2
y=32'b00000000000000000000000000111111;
x=32'b10000000000000000000000000000000;


#2
x=32'd1111111111;
y=32'd1111111111;

*/


end



always 
begin
#100 $finish;
end 


initial
begin
$monitor($time,"s=%d  a=%d  b=%d ,cout=%d   \n",s,x,y,cout1);
end
endmodule
